module add0 (a,b,q);
input a,b;
output q;
assign q = a + b;
endmodule
