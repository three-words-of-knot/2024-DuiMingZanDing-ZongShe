module full_adder(clk, ret, S, Cout, A, B, Cin);
input clk, ret;
output S;
output Cout;
input A;
input B;
input Cin;
wire A;
wire B;
wire Cin;
wire Sum1;
wire P1;
wire P2;
wire P3;
wire Cout;
wire S;
assign Sum1=A&B&Cin;
assign P1=A&B;
assign P2=B&Cin;
assign P3=A&Cin;
assign Cout=P1&P2&P3;
assign S=Sum1;
endmodule
